mstein19@remus.amherst.edu.49791:1471142699