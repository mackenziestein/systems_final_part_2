lschmidlein19@remus.amherst.edu.64055:1471142699